module displays(input modo,input decs,input segs,input resultado);
endmodule