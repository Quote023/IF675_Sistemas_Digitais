module displays(modo,decs,segs,resultado);
endmodule